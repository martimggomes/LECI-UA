library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Bin7SegDecoderDemo is
	port(SW : in std_logic_vector(3 downto 0);
			KEY : in std_logic_vector(0 downto 0);
			HEX0 : out std_logic_vector(6 downto 0));
			end Bin7SegDecoderDemo;
architecture Shell of Bin7SegDecoderDemo is
begin
Bin7SegDecoder_0: entity work.Bin7SegDecoder(Behavioral)
	port map(enable => KEY(0),
				binInput => SW,
				decOut_n => HEX0);
end Shell;				
